module Convultional_Encoder(in,out);