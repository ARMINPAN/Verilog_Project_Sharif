module Convultional_Encoder(
	
    );